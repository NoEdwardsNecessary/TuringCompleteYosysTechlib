module  \$_DFF_P_ (input D, C, output Q); DFF  _TECHMAP_REPLACE_ (.D(D), .Q(Q), .C(C), .E(1)); wire _TECHMAP_REMOVEINIT_Q_ = 1; endmodule
module  \$_DFFE_PP_ (input D, C, E, output Q); DFF  _TECHMAP_REPLACE_ (.D(D), .Q(Q), .C(C), .E(E)); wire _TECHMAP_REMOVEINIT_Q_ = 1; endmodule
